// Note: The license below is based on the template at:
// http://opensource.org/licenses/BSD-3-Clause
// Copyright (C) 2020 Regents of the University of Texas
//All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are
// met:

// o Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.

// o Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.

// o Neither the name of the copyright holders nor the names of its
//   contributors may be used to endorse or promote products derived
//   from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

// Original Author(s):
// Mertcan Temel         <mert@utexas.edu>

// DO NOT REMOVE:
// This file is generated by Temel's multiplier generator. Download from https://github.com/temelmertcan/multgen.

// Specification module to help understand what the design implements.
module U2x2 (
        input logic [1:0] IN1,
        input logic [1:0] IN2,
        input logic [0:0] IN3, //redundant

        output logic [3:0] design_res
      );
    

    WT_UB4_KS_2x2_noX mult(IN1, IN2, design_res);

    
endmodule



module WT_UB4_KS_2x2_noX(
        input logic [1:0] IN1,
        input logic [1:0] IN2,
        output logic [3:0] result);
    
    
// Creating Partial Products 

    wire [2:0] mult = {1'b0, IN1};
    wire [2:0] mcand = {1'b0, IN2};
    wire [3:0] mcand_1x;
    wire [3:0] mcand_2x;
    assign mcand_1x = {{1{mcand[2]}},  mcand};
    assign mcand_2x = {{0{mcand[2]}},  mcand, 1'b0};
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[1] mult[0] 1'b0
    wire logic select_0_0, select_e_0, select_2x_0, tcomp0, select_ne_0, select_n2x_0;
    assign select_0_0 =  &{mult[1], mult[0], 1'b0} | ~|{mult[1], mult[0], 1'b0};
    assign select_e_0 = ((~ mult[1]) & (mult[0] ^ 1'b0));
    assign select_ne_0 = mult[1] &  (mult[0] ^ 1'b0);
    assign select_2x_0 = (~ mult[1]) & mult[0] & 1'b0;
    assign select_n2x_0 = mult[1] & (~ mult[0]) & (~ 1'b0);
    reg [3:0] pp_0;
    always @(*) begin
       case (1'b1)
          select_0_0   : pp_0 = 0; 
          select_e_0   : pp_0 = mcand_1x; 
          select_2x_0  : pp_0 = mcand_2x; 
          select_n2x_0 : pp_0 = (~ mcand_2x); 
          select_ne_0  : pp_0 = (~ mcand_1x); 
          default  : pp_0 = 0; 
       endcase 
       pp_0[3] = ~pp_0[3]; // flip the MSB 
    end
    assign tcomp0 =  select_n2x_0 | select_ne_0;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[2] mult[2] mult[1]
    wire logic select_0_1, select_e_1, select_2x_1, tcomp1, select_ne_1, select_n2x_1;
    assign select_0_1 =  &{mult[2], mult[2], mult[1]} | ~|{mult[2], mult[2], mult[1]};
    assign select_e_1 = ((~ mult[2]) & (mult[2] ^ mult[1]));
    assign select_ne_1 = mult[2] &  (mult[2] ^ mult[1]);
    assign select_2x_1 = (~ mult[2]) & mult[2] & mult[1];
    assign select_n2x_1 = mult[2] & (~ mult[2]) & (~ mult[1]);
    reg [3:0] pp_1;
    always @(*) begin
       case (1'b1)
          select_0_1   : pp_1 = 0; 
          select_e_1   : pp_1 = mcand_1x; 
          select_2x_1  : pp_1 = mcand_2x; 
          select_n2x_1 : pp_1 = (~ mcand_2x); 
          select_ne_1  : pp_1 = (~ mcand_1x); 
          default  : pp_1 = 0; 
       endcase 
       pp_1[3] = ~pp_1[3]; // flip the MSB 
    end
    assign tcomp1 =  select_n2x_1 | select_ne_1;
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // pp_0[0] pp_0[1] pp_0[2] pp_0[3]   --      --    
     //   --      --    pp_1[0] pp_1[1] pp_1[2] pp_1[3] 
     // tcomp0    --    tcomp1    --      --      --    
     //   --      --      --    1'b1    1'b1      --    
    
// Creating Summation Tree 

    
    // Wallace Summation Stage 1
    logic s0 ,c0;
    ha ha0 (pp_0[0], tcomp0, s0, c0);
    logic s1 ,c1; 
    fa fa1 (pp_0[2], pp_1[0], tcomp1, s1, c1);
    logic s2 ,c2; 
    fa fa2 (pp_0[3], pp_1[1], 1'b1, s2, c2);
    
    assign result[0] = s0;
    logic [3:0] adder_result;
    KS_3 final_adder ({c1, s1, pp_0[1] }, {s2, 1'b0, c0 }, adder_result );
    assign result[3:1] = adder_result[2:0];
endmodule



module KS_3 ( 
        input logic [2:0] IN1,
        input logic [2:0] IN2,
        output logic [3:0] OUT);
    
    wire logic [2:0] p_0;
    wire logic [2:0] g_0;
    assign g_0 = IN1 & IN2;
    assign p_0 = IN1 ^ IN2;
    
// Kogge-Stone Adder 

    
    // KS stage 1
    wire logic p_1_1;
    wire logic g_1_1;
    assign p_1_1 = p_0[1] & p_0[0];
    assign g_1_1 = (p_0[1] & g_0[0]) | g_0[1];
    wire logic p_1_2;
    wire logic g_1_2;
    assign p_1_2 = p_0[2] & p_0[1];
    assign g_1_2 = (p_0[2] & g_0[1]) | g_0[2];
    
    // KS stage 2
    wire logic p_2_2;
    wire logic g_2_2;
    assign p_2_2 = p_1_2 & p_0[0];
    assign g_2_2 = (p_1_2 & g_0[0]) | g_1_2;
    
    // KS postprocess 
    assign OUT[0] = p_0[0];
    assign OUT[1] = p_0[1] ^ g_0[0];
    assign OUT[2] = p_0[2] ^ g_1_1;
    assign OUT[3] = g_2_2;
endmodule

module KS_3_spec (
        input logic [2:0] IN1,
        input logic [2:0] IN2,
        output logic adder_correct,
        output logic [3:0] spec_res);
    
    assign spec_res = IN1 + IN2;
    wire [3:0] adder_res;
    KS_3 adder(IN1, IN2, adder_res);
    assign adder_correct = ((spec_res == adder_res) ? 1 : 0);
    
endmodule



module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
endmodule

module Four2Two 
        #(parameter WIDTH=1) (
        input logic [WIDTH-1:0] in1,
        input logic [WIDTH-1:0] in2,
        input logic [WIDTH-1:0] in3,
        input logic [WIDTH-1:0] in4,
        input logic cin,
        output logic [WIDTH-1:0] sum,
        output logic [WIDTH-1:0] carry,
        output logic cout);
    
    wire logic [WIDTH:0] temp1;
    assign temp1 = {((in1 ^ in2)&in3 | in1 & ~(in1^in2)),cin};
    assign sum = ((in1 ^ in2) ^ in3 ^ in4) ^ temp1[WIDTH-1:0];
    assign carry = ((in1 ^ in2) ^ in3 ^ in4) & temp1[WIDTH-1:0] | in4 & ~((in1 ^ in2) ^ in3 ^ in4);
    assign cout = temp1[WIDTH];
endmodule




